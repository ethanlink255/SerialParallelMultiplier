magic
tech scmos
timestamp 1667532034
<< nwell >>
rect -9 48 26 105
<< ntransistor >>
rect 7 6 9 26
<< ptransistor >>
rect 7 54 9 94
<< ndiffusion >>
rect 6 6 7 26
rect 9 6 10 26
<< pdiffusion >>
rect 6 54 7 94
rect 9 54 10 94
<< ndcontact >>
rect 2 6 6 26
rect 10 6 14 26
<< pdcontact >>
rect 2 54 6 94
rect 10 54 14 94
<< psubstratepcontact >>
rect -2 -2 2 2
<< nsubstratencontact >>
rect -2 98 2 102
<< polysilicon >>
rect 7 94 9 96
rect 7 33 9 54
rect 6 29 9 33
rect 7 26 9 29
rect 7 4 9 6
<< polycontact >>
rect 2 29 6 33
<< metal1 >>
rect -2 102 18 103
rect 2 98 18 102
rect -2 97 18 98
rect 2 94 6 97
rect 2 33 6 37
rect 10 26 14 54
rect 2 3 6 6
rect -2 2 18 3
rect 2 -2 18 2
rect -2 -3 18 -2
<< m1p >>
rect 10 43 14 47
rect 2 33 6 37
<< end >>
